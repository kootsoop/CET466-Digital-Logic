/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   ���������� 4��-2�߱�����  ���ȱ�����
********************************************************************/

module my_encode(I,Y);
input [3:0] I;   ////����      �����ɿ��ؾ�����0�����£�1��δ����
output[1:0] Y;//���

reg [1:0] Y;
always@(I) //һ��I�仯��ִ��
begin             //begin end;        case endcase
	casex(I)   //���ȱ�������Ҫ��casex������  
	4'b0001:  Y=2'b00;  //I[0]Ϊ1��ʱ�����Ϊ0
	4'b001x:  Y=2'b01;  //I[1]Ϊ1��ʱ�����Ϊ1
	4'b01xx:  Y=2'b10; //I[2]Ϊ1��ʱ�����Ϊ2
	4'b1xxx:  Y=2'b11;//I[3]Ϊ1��ʱ�����Ϊ3
     default:   Y=2'b00; //����״̬�Ĵ���
  endcase
end	
endmodule
