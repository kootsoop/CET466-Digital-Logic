/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.07
**�汾�ţ�     version 1.0
**����������   led����˸ʵ�飬4��LED�ƻ���һ��Ƶ����˸
********************************************************************/




module led_twinkle(led,clk);// ģ�������˿ڲ���
	output [3:0] led;
	input clk;
	reg[3:0] led;// ����˿ڶ���Ϊ�Ĵ�����
	reg[24:0] counter;  // �м����counter����Ϊ�Ĵ�����
	
	always@(posedge clk)//��ʱ�Ӹ�������
		begin // ˳����䣬��endֹ
			counter<=counter+1;  //<=�� =����
		    //if(counter==25'b1011111010111100001000000) //�б�counter�е���ֵΪ25000000ʱ
		    if(counter==25'd25000000)
			
				begin	
					led<=~led;// led[0]-led[3]��תһ��
			 		counter<=0;//���¼���
				end   
		end
endmodule
	