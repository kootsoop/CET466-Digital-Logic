altpll0_inst : altpll0 PORT MAP (
		inclk0	 => inclk0_sig,
		c1	 => c1_sig,
		c2	 => c2_sig
	);
