/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������    ȫ������������������������Ӷ���	     
********************************************************************/

module full_adder(
    A,						//����ѡ���ַ�ɿ��ؾ�����0�����£�1��δ����
	B,						//����ѡ���ַ�ɿ��ؾ�����0�����£�1��δ����
	Ci,						//��λ��λֵ����ѡ���ַ�ɿ��ؾ�����0�����£�1��δ����
	
	S,						//��λ�ͣ������0��������1��Ϩ��
	Co						//���λ��λ�������0��������1��Ϩ��
    );
input			A;				//����˿�
input			B;				//����˿�
input			Ci;				//����˿�

output		S;				//����˿�
output		Co;				//����˿�

wire			C0;				//����˵��
wire			C1;				//����˵��

assign Co = C0 | C1;				//���ţ������������������ȫ�������

half_adder half_adder_0(			//��һ�����������
	.A(A),					//�˿�A
	.B(B),					//�˿�B
	
	.S(A0),					//�˿�S
	.C(C0)					//�˿�C
	);
	
half_adder half_adder_1(
	.A(A0),					//�˿�A	
	.B(Ci),					//�˿�B
	
	.S(S),						//�˿�S			
	.C(C1)					//�˿�C	
	);

endmodule
