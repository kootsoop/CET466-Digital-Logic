/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   ���뿪����������LED  
������뿪������ȥ1,��ô����LED1
������뿪������ȥ2,��ô����LED2
********************************************************************/


module ckey_led(ckey,LED);
  input  [4:1] ckey;                   // ckey[1]  ~ ckey[4]
  output [4:1] LED;                    // LED[1] ~ LED[4]
   

// ��������LED[1]����LED[4]���ң���1����0��
// ��������ckey��Ϊ0���ر�Ϊ1
assign LED = ckey;

endmodule